module IntXbar(
  output logic [2:0] o,
  input logic i);
endmodule
